module main
import os
// import fs

fn main() {
	os.execute("")
	
}