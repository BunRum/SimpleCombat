module main
import os
// import fs

fn rec(dir) {
	f := {[]}
	
	files := os.glob() or {[]}
}

fn main() {
	files := os.glob() or {[]}
	print(files)
	// os.glob()
}