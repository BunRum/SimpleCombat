module main

fn main() {
	print("how amazing")
}