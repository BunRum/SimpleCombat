module main
import os
// import fs

fn rec(dir) {
	f := 
}

fn main() {
	files := os.glob() or {[]}
	print(files)
	// os.glob()
}