module main
import os
// import fs

fn rec(dir) {
	
}

fn main() {
	files := os.glob() or {[]}
	print(files)
	// os.glob()
}