module main
import os

fn main() {
	os.execute("")
}