module main
import os
// import fs

fn main() {
	print(os.dir("./"))
}