module main
import os
// import fs

fn rec(dir) {
	f := {[]}
	for
}

fn main() {
	files := os.glob() or {[]}
	print(files)
	// os.glob()
}